module fixedtofloat
(
	clk,
	clken,
	fixedin,
	floatout
);

	input clk;
	input	clken;
	input signed [27:0] fixedin;
	output reg [31:0] floatout;
	reg [27:0] internal;
	reg sign;
	
	
	
	always @ (posedge clk) 	begin
		if(fixedin[27]) begin
			internal <= ~fixedin + 1;
			sign <= 1'b1;
		end
		else begin
			internal <= fixedin;
			sign <= 1'b0;
		end
			
		case(fixedin)
			28'b01xxxxxxxxxxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd127, internal[25:3] };
			end
			28'b001xxxxxxxxxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd126, internal[24:2]};
			end
			28'b0001xxxxxxxxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd125, internal[23:1]};
			end
			28'b00001xxxxxxxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd124, internal[22:0]};
			end
			28'b000001xxxxxxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd123, internal[21:0], 1'b0};
			end
			28'b0000001xxxxxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd122, internal[20:0], 2'b0};
			end
			28'b00000001xxxxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd121, internal[19:0], 3'b0};
			end
			28'b000000001xxxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd120, internal[18:0], 4'b0};
			end
			28'b0000000001xxxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd119, internal[17:0], 5'b0};
			end
			28'b00000000001xxxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd118, internal[16:0], 6'b0};
			end  
			28'b000000000001xxxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd117, internal[15:0], 7'b0};
			end
			28'b0000000000001xxxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd116, internal[14:0], 8'b0};
			end
			28'b00000000000001xxxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd115, internal[13:0], 9'b0};
			end
			28'b000000000000001xxxxxxxxxxxxx: begin
				floatout <= {sign, 8'd114, internal[12:0], 10'b0};
			end
			28'b0000000000000001xxxxxxxxxxxx: begin
				floatout <= {sign, 8'd113, internal[11:0], 11'b0};
			end
			28'b00000000000000001xxxxxxxxxxx: begin
				floatout <= {sign, 8'd112, internal[10:0], 12'b0};
			end
			28'b000000000000000001xxxxxxxxxx: begin
				floatout <= {sign, 8'd111, internal[9:0], 13'b0};
			end
			28'b0000000000000000001xxxxxxxxx: begin
				floatout <= {sign, 8'd110, internal[8:0], 14'b0};
			end
			28'b00000000000000000001xxxxxxxx: begin
				floatout <= {sign, 8'd109, internal[7:0], 15'b0};
			end
			28'b000000000000000000001xxxxxxx: begin
				floatout <= {sign, 8'd108, internal[6:0], 16'b0};
			end
			28'b0000000000000000000001xxxxxx: begin
				floatout <= {sign, 8'd107, internal[5:0], 17'b0};
			end
			28'b00000000000000000000001xxxxx: begin
				floatout <= {sign, 8'd106, internal[4:0], 18'b0};
			end
			28'b000000000000000000000001xxxx: begin
				floatout <= {sign, 8'd105, internal[3:0], 19'b0};
			end
			28'b0000000000000000000000001xxx: begin
				floatout <= {sign, 8'd104, internal[2:0], 20'b0};
			end
			28'b00000000000000000000000001xx: begin
				floatout <= {sign, 8'd103, internal[1:0], 21'b0};
			end
			28'b000000000000000000000000001x: begin
				floatout <= {sign, 8'd102, internal[0], 22'b0};
			end
			28'b0000000000000000000000000001: begin
				floatout <= {sign, 8'd101, 23'd0};
			end
			28'b0000000000000000000000000000: begin
				floatout <= {sign, 8'd0, 23'd0};
			end
	endcase
	
	
	end
endmodule

/*


0d58fa94 goes to
3f558fa9

001101010110001111101010010100
00111111010101011000111110101001
SeeeeeeeeMMMMMMMMMMMMMMMMMMMMMMM


001101010110001111101010010100

=> 10101011000111110101001 */ 